

`define N_TESTS 100000
module division_tb;
	reg [31:0] a_operand;
	reg [31:0] b_operand;
	reg        En;
	wire [31:0] result;


	FPU_MUL DUT(.En(En),.Rs1(a_operand),.Rs2(b_operand));

	initial  
	begin 
			En   = 1'b1;

			a_operand =  32'b01000011100011110110000000000000;
			b_operand =  32'b10111111100100101000000000000000;
				
			#1
			
			a_operand = 32'b11000001011000000000000000000000;
			b_operand =  32'b11000000000000000000000000000000;
			
			
					
			#1

			
			a_operand = 32'b01000000010000000000000000000000;
			b_operand =  32'b01000000000000000000000000000000;
			
			#1

			
			a_operand = 32'b11000001100101000000000000000000;
			b_operand = 32'b01000000000000000000000000000000;
			
			#1
	
			
			a_operand = 32'b01000001101100000000000000000000;
			b_operand =  32'b01000000111000000000000000000000;
			
			#1

			
			a_operand = 32'b01000000001100000000000000000000;
			b_operand =  32'b01000000110010110101110000101001;
			
		#1

			
			a_operand = 32'b01000010111111100001000000000000;
			b_operand =  32'b01000001100001111000000000000000;
			
			#1

			
			a_operand = 32'b01000010100011111100000000000000;
			b_operand =  32'b01000000110010000000000000000000;
			
			#1


	$stop;
	end 




endmodule